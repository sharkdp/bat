[38;2;190;132;255m`timescale[0m[38;2;248;248;242m [0m[38;2;190;132;255m1ns[0m[38;2;249;38;114m/[0m[38;2;190;132;255m1ps[0m

[38;2;117;113;94m//[0m[38;2;117;113;94m Design Code[0m
[38;2;249;38;114mmodule[0m[38;2;248;248;242m [0m[38;2;166;226;46mADDER[0m[38;2;248;248;242m([0m
[3;38;2;166;226;46m    input[0m[38;2;248;248;242m clk,[0m
[3;38;2;166;226;46m    input[0m[38;2;248;248;242m [[0m[38;2;190;132;255m7[0m[38;2;249;38;114m:[0m[38;2;190;132;255m0[0m[38;2;248;248;242m]	a,[0m
[3;38;2;166;226;46m    input[0m[38;2;248;248;242m [[0m[38;2;190;132;255m7[0m[38;2;249;38;114m:[0m[38;2;190;132;255m0[0m[38;2;248;248;242m]	b,[0m
[3;38;2;166;226;46m    input[0m[38;2;248;248;242m bIsPos,[0m
[38;2;248;248;242m    [0m[3;38;2;166;226;46moutput[0m[38;2;248;248;242m [0m[3;38;2;102;217;239mreg[0m[38;2;248;248;242m [[0m[38;2;190;132;255m8[0m[38;2;249;38;114m:[0m[38;2;190;132;255m0[0m[38;2;248;248;242m] result[0m
[38;2;248;248;242m);[0m

[38;2;248;248;242m    [0m[38;2;249;38;114malways[0m[38;2;248;248;242m [0m[38;2;249;38;114m@[0m[38;2;248;248;242m ([0m[38;2;249;38;114mposedge[0m[38;2;248;248;242m clk) [0m[38;2;249;38;114mbegin[0m
[38;2;248;248;242m        [0m[38;2;249;38;114mif[0m[38;2;248;248;242m (bIsPos) [0m[38;2;249;38;114mbegin[0m[38;2;248;248;242m	[0m
[38;2;248;248;242m            result [0m[38;2;249;38;114m<=[0m[38;2;248;248;242m a [0m[38;2;249;38;114m+[0m[38;2;248;248;242m b;[0m
[38;2;248;248;242m        [0m[38;2;249;38;114mend[0m[38;2;248;248;242m [0m[38;2;249;38;114melse[0m[38;2;248;248;242m [0m[38;2;249;38;114mbegin[0m
[38;2;248;248;242m            result [0m[38;2;249;38;114m<=[0m[38;2;248;248;242m a [0m[38;2;249;38;114m-[0m[38;2;248;248;242m b;[0m
[38;2;248;248;242m        [0m[38;2;249;38;114mend[0m
[38;2;248;248;242m    [0m[38;2;249;38;114mend[0m

[38;2;249;38;114mendmodule[0m[38;2;249;38;114m:[0m[38;2;248;248;242m [0m[38;2;166;226;46mADDER[0m

[38;2;249;38;114minterface[0m[38;2;248;248;242m [0m[38;2;166;226;46madder_if[0m[38;2;248;248;242m([0m
[38;2;248;248;242m    [0m[3;38;2;166;226;46minput[0m[38;2;248;248;242m [0m[3;38;2;102;217;239mbit[0m[38;2;248;248;242m clk,[0m
[3;38;2;166;226;46m    input[0m[38;2;248;248;242m [[0m[38;2;190;132;255m7[0m[38;2;249;38;114m:[0m[38;2;190;132;255m0[0m[38;2;248;248;242m] a,[0m
[3;38;2;166;226;46m    input[0m[38;2;248;248;242m [[0m[38;2;190;132;255m7[0m[38;2;249;38;114m:[0m[38;2;190;132;255m0[0m[38;2;248;248;242m] b,[0m
[3;38;2;166;226;46m    input[0m[38;2;248;248;242m bIsPos,[0m
[3;38;2;166;226;46m    input[0m[38;2;248;248;242m [[0m[38;2;190;132;255m8[0m[38;2;249;38;114m:[0m[38;2;190;132;255m0[0m[38;2;248;248;242m] result[0m
[38;2;248;248;242m);[0m

[38;2;248;248;242m    [0m[38;2;249;38;114mclocking[0m[38;2;248;248;242m cb [0m[38;2;249;38;114m@[0m[38;2;248;248;242m([0m[38;2;249;38;114mposedge[0m[38;2;248;248;242m clk);[0m
[3;38;2;166;226;46m        output[0m[38;2;248;248;242m a;[0m
[3;38;2;166;226;46m        output[0m[38;2;248;248;242m b;[0m
[3;38;2;166;226;46m        output[0m[38;2;248;248;242m bIsPos;[0m
[3;38;2;166;226;46m        input[0m[38;2;248;248;242m result;[0m
[38;2;248;248;242m    [0m[38;2;249;38;114mendclocking[0m[38;2;248;248;242m [0m[38;2;249;38;114m:[0m[38;2;248;248;242m [0m[38;2;166;226;46mcb[0m

[38;2;249;38;114mendinterface[0m[38;2;249;38;114m:[0m[38;2;248;248;242m [0m[38;2;166;226;46madder_if[0m


[38;2;249;38;114mbind[0m[38;2;248;248;242m ADDER [0m[3;38;2;102;217;239madder_if[0m[38;2;248;248;242m [0m[38;2;166;226;46mmy_adder_if[0m[38;2;248;248;242m([0m
[38;2;248;248;242m    .[0m[38;2;102;217;239mclk[0m[38;2;248;248;242m(clk),[0m
[38;2;248;248;242m    .[0m[38;2;102;217;239ma[0m[38;2;248;248;242m(a),[0m
[38;2;248;248;242m    .[0m[38;2;102;217;239mb[0m[38;2;248;248;242m(b),[0m
[38;2;248;248;242m    .[0m[38;2;102;217;239mbIsPos[0m[38;2;248;248;242m(bIsPos),[0m
[38;2;248;248;242m    .[0m[38;2;102;217;239mresult[0m[38;2;248;248;242m(result)[0m
[38;2;248;248;242m);[0m


[38;2;117;113;94m//[0m[38;2;117;113;94m Testbench Code[0m
[38;2;249;38;114mimport[0m[38;2;248;248;242m [0m[3;38;2;166;226;46muvm_pkg[0m[38;2;249;38;114m::[0m[38;2;249;38;114m*[0m[38;2;248;248;242m;[0m
[38;2;190;132;255m`include[0m[38;2;248;248;242m [0m[38;2;230;219;116m"[0m[38;2;230;219;116muvm_macros.svh[0m[38;2;230;219;116m"[0m

[38;2;249;38;114mclass[0m[38;2;248;248;242m [0m[38;2;166;226;46mtestbench_env[0m[38;2;248;248;242m [0m[38;2;249;38;114mextends[0m[38;2;248;248;242m [0m[3;4;38;2;166;226;46muvm_env[0m[38;2;248;248;242m;[0m

[38;2;248;248;242m    [0m[38;2;249;38;114mvirtual [0m[3;38;2;102;217;239madder_if[0m[38;2;248;248;242m [0m[38;2;248;248;242mm_if;[0m

[38;2;248;248;242m    [0m[38;2;249;38;114mfunction[0m[38;2;248;248;242m [0m[38;2;166;226;46mnew[0m[38;2;248;248;242m([0m[3;38;2;102;217;239mstring[0m[38;2;248;248;242m name, [0m[3;38;2;102;217;239muvm_component[0m[38;2;248;248;242m parent [0m[38;2;249;38;114m=[0m[38;2;248;248;242m [0m[38;2;102;217;239mnull[0m[38;2;248;248;242m)[0m[38;2;248;248;242m;[0m
[38;2;248;248;242m        [0m[38;2;249;38;114msuper[0m[38;2;248;248;242m.[0m[38;2;249;38;114mnew[0m[38;2;248;248;242m(name, parent);[0m
[38;2;248;248;242m    [0m[38;2;249;38;114mendfunction[0m
[38;2;248;248;242m    [0m
[38;2;248;248;242m    [0m[38;2;249;38;114mfunction[0m[3;38;2;102;217;239m void[0m[38;2;248;248;242m [0m[38;2;166;226;46mconnect_phase[0m[38;2;248;248;242m([0m[3;38;2;102;217;239muvm_phase[0m[38;2;248;248;242m phase[0m[38;2;248;248;242m)[0m[38;2;248;248;242m;[0m
[38;2;248;248;242m        [0m[38;2;249;38;114massert[0m[38;2;248;248;242m(uvm_resource_db[0m[38;2;249;38;114m#[0m[38;2;248;248;242m([0m[38;2;249;38;114mvirtual[0m[38;2;248;248;242m adder_if)[0m[38;2;249;38;114m:[0m[38;2;249;38;114m:[0m[38;2;102;217;239mread_by_name[0m[38;2;248;248;242m([0m[38;2;102;217;239mget_full_name[0m[38;2;248;248;242m(), [0m[38;2;230;219;116m"[0m[38;2;230;219;116madder_if[0m[38;2;230;219;116m"[0m[38;2;248;248;242m, m_if));[0m
[38;2;248;248;242m    [0m[38;2;249;38;114mendfunction[0m[38;2;249;38;114m:[0m[38;2;248;248;242m [0m[38;2;166;226;46mconnect_phase[0m

[38;2;248;248;242m    [0m[38;2;249;38;114mtask[0m[38;2;248;248;242m [0m[38;2;166;226;46mrun_phase[0m[38;2;248;248;242m([0m[3;38;2;102;217;239muvm_phase[0m[38;2;248;248;242m phase[0m[38;2;248;248;242m)[0m[38;2;248;248;242m;[0m
[38;2;248;248;242m        phase.[0m[38;2;102;217;239mraise_objection[0m[38;2;248;248;242m([0m[38;2;249;38;114mthis[0m[38;2;248;248;242m);[0m
[38;2;248;248;242m        [0m[38;2;190;132;255m`uvm_info[0m[38;2;248;248;242m([0m[38;2;102;217;239mget_name[0m[38;2;248;248;242m(), [0m[38;2;230;219;116m"[0m[38;2;230;219;116mStarting test![0m[38;2;230;219;116m"[0m[38;2;248;248;242m, [0m[38;2;190;132;255mUVM_HIGH[0m[38;2;248;248;242m);[0m
[38;2;248;248;242m        [0m[38;2;249;38;114mbegin[0m
[3;38;2;102;217;239m            int[0m[38;2;248;248;242m a [0m[38;2;249;38;114m=[0m[38;2;248;248;242m [0m[38;2;190;132;255m8'h4[0m[38;2;248;248;242m, b [0m[38;2;249;38;114m=[0m[38;2;248;248;242m [0m[38;2;190;132;255m8'h5[0m[38;2;248;248;242m;[0m
[38;2;248;248;242m            [0m[38;2;249;38;114m@[0m[38;2;248;248;242m(m_if.cb);[0m
[38;2;248;248;242m            m_if.cb.a [0m[38;2;249;38;114m<=[0m[38;2;248;248;242m a;[0m
[38;2;248;248;242m            m_if.cb.b [0m[38;2;249;38;114m<=[0m[38;2;248;248;242m b;[0m
[38;2;248;248;242m            m_if.cb.bIsPos [0m[38;2;249;38;114m<=[0m[38;2;248;248;242m [0m[38;2;190;132;255m1'b1[0m[38;2;248;248;242m;[0m
[38;2;248;248;242m            [0m[38;2;249;38;114mrepeat[0m[38;2;248;248;242m([0m[38;2;190;132;255m2[0m[38;2;248;248;242m) [0m[38;2;249;38;114m@[0m[38;2;248;248;242m(m_if.cb);[0m
[38;2;248;248;242m            [0m[38;2;190;132;255m`uvm_info[0m[38;2;248;248;242m([0m[38;2;102;217;239mget_name[0m[38;2;248;248;242m(), [0m[38;2;102;217;239m$sformatf[0m[38;2;248;248;242m([0m[38;2;230;219;116m"[0m[38;2;190;132;255m%0d[0m[38;2;230;219;116m + [0m[38;2;190;132;255m%0d[0m[38;2;230;219;116m = [0m[38;2;190;132;255m%0d[0m[38;2;230;219;116m"[0m[38;2;248;248;242m, a, b, m_if.cb.result), [0m[38;2;190;132;255mUVM_LOW[0m[38;2;248;248;242m);[0m
[38;2;248;248;242m        [0m[38;2;249;38;114mend[0m
[38;2;248;248;242m        [0m[38;2;190;132;255m`uvm_info[0m[38;2;248;248;242m([0m[38;2;102;217;239mget_name[0m[38;2;248;248;242m(), [0m[38;2;230;219;116m"[0m[38;2;230;219;116mEnding test![0m[38;2;230;219;116m"[0m[38;2;248;248;242m, [0m[38;2;190;132;255mUVM_HIGH[0m[38;2;248;248;242m);[0m
[38;2;248;248;242m        phase.[0m[38;2;102;217;239mdrop_objection[0m[38;2;248;248;242m([0m[38;2;249;38;114mthis[0m[38;2;248;248;242m);[0m
[38;2;248;248;242m    [0m[38;2;249;38;114mendtask[0m[38;2;249;38;114m:[0m[38;2;248;248;242m [0m[38;2;166;226;46mrun_phase[0m
[38;2;249;38;114mendclass[0m


[38;2;249;38;114mmodule[0m[38;2;248;248;242m [0m[38;2;166;226;46mtop[0m[38;2;248;248;242m;[0m

[3;38;2;102;217;239m    bit[0m[38;2;248;248;242m clk;[0m
[38;2;248;248;242m    [0m[3;38;2;102;217;239menv[0m[38;2;248;248;242m [0m[38;2;248;248;242menvironment;[0m
[38;2;248;248;242m    [0m[3;38;2;102;217;239mADDER[0m[38;2;248;248;242m [0m[38;2;166;226;46mdut[0m[38;2;248;248;242m(.[0m[38;2;102;217;239mclk[0m[38;2;248;248;242m (clk));[0m

[38;2;248;248;242m    [0m[38;2;249;38;114minitial[0m[38;2;248;248;242m [0m[38;2;249;38;114mbegin[0m
[38;2;248;248;242m        [0m[38;2;248;248;242menvironment [0m[38;2;249;38;114m=[0m[38;2;248;248;242m [0m[38;2;249;38;114mnew[0m[38;2;248;248;242m([0m[38;2;230;219;116m"[0m[38;2;230;219;116mtestbench_env[0m[38;2;230;219;116m"[0m[38;2;248;248;242m);[0m
[38;2;248;248;242m        [0m[3;38;2;102;217;239muvm_resource_db[0m[38;2;249;38;114m#[0m[38;2;248;248;242m([0m[38;2;249;38;114mvirtual[0m[38;2;248;248;242m adder_if)[0m[38;2;249;38;114m:[0m[38;2;249;38;114m:[0m[38;2;102;217;239mset[0m[38;2;248;248;242m([0m[38;2;230;219;116m"[0m[38;2;230;219;116menv[0m[38;2;230;219;116m"[0m[38;2;248;248;242m, [0m[38;2;230;219;116m"[0m[38;2;230;219;116madder_if[0m[38;2;230;219;116m"[0m[38;2;248;248;242m, dut.my_adder_if);[0m
[38;2;248;248;242m        [0m[38;2;248;248;242mclk [0m[38;2;249;38;114m=[0m[38;2;248;248;242m [0m[38;2;190;132;255m0[0m[38;2;248;248;242m;[0m
[38;2;248;248;242m        [0m[38;2;102;217;239mrun_test[0m[38;2;248;248;242m();[0m
[38;2;248;248;242m    [0m[38;2;249;38;114mend[0m

[38;2;248;248;242m    [0m[38;2;117;113;94m//[0m[38;2;117;113;94m Clock generation	[0m
[38;2;248;248;242m    [0m[38;2;249;38;114minitial[0m[38;2;248;248;242m [0m[38;2;249;38;114mbegin[0m
[38;2;248;248;242m        [0m[38;2;249;38;114mforever[0m[38;2;248;248;242m [0m[38;2;249;38;114mbegin[0m
[38;2;248;248;242m            [0m[38;2;249;38;114m#[0m[38;2;248;248;242m([0m[38;2;190;132;255m1[0m[38;2;248;248;242m) clk [0m[38;2;249;38;114m=[0m[38;2;248;248;242m [0m[38;2;249;38;114m~[0m[38;2;248;248;242mclk;[0m
[38;2;248;248;242m        [0m[38;2;249;38;114mend[0m
[38;2;248;248;242m    [0m[38;2;249;38;114mend[0m
[38;2;248;248;242m    [0m
[38;2;249;38;114mendmodule[0m
