[38;2;117;113;94m--[0m[38;2;117;113;94m This is a single-line comment[0m

[38;2;249;38;114mlibrary[0m[38;2;248;248;242m [0m[38;2;248;248;242mIEEE[0m[38;2;248;248;242m;[0m
[38;2;249;38;114muse[0m[38;2;248;248;242m [0m[38;2;248;248;242mIEEE[0m[38;2;248;248;242m.[0m[38;2;248;248;242mSTD_LOGIC_1164[0m[38;2;248;248;242m.[0m[38;2;249;38;114mALL[0m[38;2;248;248;242m;[0m
[38;2;249;38;114muse[0m[38;2;248;248;242m [0m[38;2;248;248;242mIEEE[0m[38;2;248;248;242m.[0m[38;2;248;248;242mNUMERIC_STD[0m[38;2;248;248;242m.[0m[38;2;249;38;114mALL[0m[38;2;248;248;242m;[0m

[38;2;249;38;114mentity[0m[38;2;248;248;242m [0m[38;2;166;226;46mSyntaxTest[0m[38;2;248;248;242m [0m[38;2;249;38;114mis[0m
[38;2;248;248;242m    [0m[38;2;249;38;114mgeneric[0m[38;2;248;248;242m [0m[38;2;248;248;242m([0m
[38;2;248;248;242m        [0m[38;2;248;248;242mDATA_WIDTH [0m[38;2;248;248;242m:[0m[38;2;248;248;242m [0m[3;38;2;102;217;239minteger[0m[38;2;248;248;242m [0m[38;2;249;38;114m:=[0m[38;2;248;248;242m [0m[38;2;190;132;255m8[0m
[38;2;248;248;242m    [0m[38;2;248;248;242m)[0m[38;2;248;248;242m;[0m
[38;2;248;248;242m    [0m[38;2;249;38;114mport[0m[38;2;248;248;242m [0m[38;2;248;248;242m([0m
[38;2;248;248;242m        [0m[38;2;248;248;242mclk     [0m[38;2;248;248;242m:[0m[38;2;248;248;242m [0m[38;2;249;38;114min[0m[38;2;248;248;242m  [0m[3;38;2;102;217;239mstd_logic[0m[38;2;248;248;242m;[0m
[38;2;248;248;242m        [0m[38;2;248;248;242mrst     [0m[38;2;248;248;242m:[0m[38;2;248;248;242m [0m[38;2;249;38;114min[0m[38;2;248;248;242m  [0m[3;38;2;102;217;239mstd_logic[0m[38;2;248;248;242m;[0m
[38;2;248;248;242m        [0m[38;2;248;248;242ma[0m[38;2;248;248;242m,[0m[38;2;248;248;242m [0m[38;2;248;248;242mb    [0m[38;2;248;248;242m:[0m[38;2;248;248;242m [0m[38;2;249;38;114min[0m[38;2;248;248;242m  [0m[3;38;2;102;217;239mstd_logic_vector[0m[38;2;248;248;242m([0m[38;2;248;248;242mDATA_WIDTH [0m[38;2;249;38;114m-[0m[38;2;248;248;242m [0m[38;2;190;132;255m1[0m[38;2;248;248;242m [0m[38;2;249;38;114mdownto[0m[38;2;248;248;242m [0m[38;2;190;132;255m0[0m[38;2;248;248;242m)[0m[38;2;248;248;242m;[0m
[38;2;248;248;242m        [0m[38;2;248;248;242msel     [0m[38;2;248;248;242m:[0m[38;2;248;248;242m [0m[38;2;249;38;114min[0m[38;2;248;248;242m  [0m[3;38;2;102;217;239mstd_logic[0m[38;2;248;248;242m;[0m
[38;2;248;248;242m        [0m[38;2;248;248;242mresult  [0m[38;2;248;248;242m:[0m[38;2;248;248;242m [0m[38;2;249;38;114mout[0m[38;2;248;248;242m [0m[3;38;2;102;217;239mstd_logic_vector[0m[38;2;248;248;242m([0m[38;2;248;248;242mDATA_WIDTH [0m[38;2;249;38;114m-[0m[38;2;248;248;242m [0m[38;2;190;132;255m1[0m[38;2;248;248;242m [0m[38;2;249;38;114mdownto[0m[38;2;248;248;242m [0m[38;2;190;132;255m0[0m[38;2;248;248;242m)[0m[38;2;248;248;242m;[0m
[38;2;248;248;242m        [0m[38;2;248;248;242mflag    [0m[38;2;248;248;242m:[0m[38;2;248;248;242m [0m[38;2;249;38;114mout[0m[38;2;248;248;242m [0m[3;38;2;102;217;239mstd_logic[0m
[38;2;248;248;242m    [0m[38;2;248;248;242m)[0m[38;2;248;248;242m;[0m
[38;2;249;38;114mend[0m[38;2;248;248;242m [0m[38;2;166;226;46mSyntaxTest[0m[38;2;248;248;242m;[0m

[38;2;249;38;114marchitecture[0m[38;2;248;248;242m [0m[38;2;166;226;46mBehavioral[0m[38;2;248;248;242m [0m[38;2;249;38;114mof[0m[38;2;248;248;242m [0m[38;2;166;226;46mSyntaxTest[0m[38;2;248;248;242m [0m[38;2;249;38;114mis[0m

[38;2;248;248;242m    [0m[38;2;249;38;114msignal[0m[38;2;248;248;242m tmp [0m[38;2;248;248;242m:[0m[38;2;248;248;242m [0m[3;38;2;102;217;239mstd_logic_vector[0m[38;2;248;248;242m([0m[38;2;248;248;242mDATA_WIDTH [0m[38;2;249;38;114m-[0m[38;2;248;248;242m [0m[38;2;190;132;255m1[0m[38;2;248;248;242m [0m[38;2;249;38;114mdownto[0m[38;2;248;248;242m [0m[38;2;190;132;255m0[0m[38;2;248;248;242m)[0m[38;2;248;248;242m;[0m
[38;2;248;248;242m    [0m[38;2;249;38;114msignal[0m[38;2;248;248;242m done [0m[38;2;248;248;242m:[0m[38;2;248;248;242m [0m[3;38;2;102;217;239mstd_logic[0m[38;2;248;248;242m [0m[38;2;249;38;114m:=[0m[38;2;248;248;242m [0m[38;2;190;132;255m'0'[0m[38;2;248;248;242m;[0m

[38;2;248;248;242m    [0m[38;2;249;38;114mtype[0m[38;2;248;248;242m [0m[38;2;166;226;46mstate_type[0m[38;2;248;248;242m [0m[38;2;249;38;114mis[0m[38;2;248;248;242m [0m[38;2;248;248;242m([0m[38;2;248;248;242mIDLE[0m[38;2;248;248;242m,[0m[38;2;248;248;242m LOAD[0m[38;2;248;248;242m,[0m[38;2;248;248;242m EXECUTE[0m[38;2;248;248;242m,[0m[38;2;248;248;242m DONE[0m[38;2;248;248;242m)[0m[38;2;248;248;242m;[0m
[38;2;248;248;242m    [0m[38;2;249;38;114msignal[0m[38;2;248;248;242m state [0m[38;2;248;248;242m:[0m[38;2;248;248;242m [0m[3;38;2;102;217;239mstate_type[0m[38;2;248;248;242m [0m[38;2;249;38;114m:=[0m[38;2;248;248;242m [0m[3;38;2;102;217;239mIDLE[0m[38;2;248;248;242m;[0m

[38;2;249;38;114mbegin[0m

[38;2;248;248;242m    [0m[38;2;249;38;114mprocess[0m[38;2;248;248;242m([0m[38;2;248;248;242mclk[0m[38;2;248;248;242m,[0m[38;2;248;248;242m rst[0m[38;2;248;248;242m)[0m
[38;2;248;248;242m        [0m[38;2;249;38;114mvariable[0m[38;2;248;248;242m i [0m[38;2;248;248;242m:[0m[38;2;248;248;242m [0m[3;38;2;102;217;239minteger[0m[38;2;248;248;242m [0m[38;2;249;38;114m:=[0m[38;2;248;248;242m [0m[38;2;190;132;255m0[0m[38;2;248;248;242m;[0m
[38;2;248;248;242m    [0m[38;2;249;38;114mbegin[0m
[38;2;248;248;242m        [0m[38;2;249;38;114mif[0m[38;2;248;248;242m rst [0m[38;2;249;38;114m=[0m[38;2;248;248;242m [0m[38;2;190;132;255m'1'[0m[38;2;248;248;242m [0m[38;2;249;38;114mthen[0m
[38;2;248;248;242m            tmp   [0m[38;2;249;38;114m<=[0m[38;2;248;248;242m [0m[38;2;248;248;242m([0m[38;2;249;38;114mothers[0m[38;2;248;248;242m [0m[38;2;249;38;114m=>[0m[38;2;248;248;242m [0m[38;2;190;132;255m'0'[0m[38;2;248;248;242m)[0m[38;2;248;248;242m;[0m
[38;2;248;248;242m            flag  [0m[38;2;249;38;114m<=[0m[38;2;248;248;242m [0m[38;2;190;132;255m'0'[0m[38;2;248;248;242m;[0m
[38;2;248;248;242m            state [0m[38;2;249;38;114m<=[0m[38;2;248;248;242m IDLE[0m[38;2;248;248;242m;[0m

[38;2;248;248;242m        [0m[38;2;249;38;114melsif[0m[38;2;248;248;242m [0m[38;2;102;217;239mrising_edge[0m[38;2;248;248;242m([0m[38;2;248;248;242mclk[0m[38;2;248;248;242m)[0m[38;2;248;248;242m [0m[38;2;249;38;114mthen[0m
[38;2;248;248;242m            [0m[38;2;249;38;114mcase[0m[38;2;248;248;242m state [0m[38;2;249;38;114mis[0m
[38;2;248;248;242m                [0m[38;2;249;38;114mwhen[0m[38;2;248;248;242m IDLE [0m[38;2;249;38;114m=>[0m
[38;2;248;248;242m                    [0m[38;2;249;38;114mif[0m[38;2;248;248;242m sel [0m[38;2;249;38;114m=[0m[38;2;248;248;242m [0m[38;2;190;132;255m'1'[0m[38;2;248;248;242m [0m[38;2;249;38;114mthen[0m
[38;2;248;248;242m                        tmp [0m[38;2;249;38;114m<=[0m[38;2;248;248;242m a [0m[38;2;249;38;114mand[0m[38;2;248;248;242m b[0m[38;2;248;248;242m;[0m
[38;2;248;248;242m                        state [0m[38;2;249;38;114m<=[0m[38;2;248;248;242m EXECUTE[0m[38;2;248;248;242m;[0m
[38;2;248;248;242m                    [0m[38;2;249;38;114melse[0m
[38;2;248;248;242m                        tmp [0m[38;2;249;38;114m<=[0m[38;2;248;248;242m a [0m[38;2;249;38;114mor[0m[38;2;248;248;242m b[0m[38;2;248;248;242m;[0m
[38;2;248;248;242m                        state [0m[38;2;249;38;114m<=[0m[38;2;248;248;242m LOAD[0m[38;2;248;248;242m;[0m
[38;2;248;248;242m                    [0m[38;2;249;38;114mend[0m[38;2;248;248;242m [0m[38;2;249;38;114mif[0m[38;2;248;248;242m;[0m

[38;2;248;248;242m                [0m[38;2;249;38;114mwhen[0m[38;2;248;248;242m LOAD [0m[38;2;249;38;114m=>[0m
[38;2;248;248;242m                    tmp [0m[38;2;249;38;114m<=[0m[38;2;248;248;242m a [0m[38;2;249;38;114mxor[0m[38;2;248;248;242m b[0m[38;2;248;248;242m;[0m
[38;2;248;248;242m                    state [0m[38;2;249;38;114m<=[0m[38;2;248;248;242m EXECUTE[0m[38;2;248;248;242m;[0m

[38;2;248;248;242m                [0m[38;2;249;38;114mwhen[0m[38;2;248;248;242m EXECUTE [0m[38;2;249;38;114m=>[0m
[38;2;248;248;242m                    [0m[38;2;249;38;114mif[0m[38;2;248;248;242m i [0m[38;2;249;38;114m<[0m[38;2;248;248;242m DATA_WIDTH [0m[38;2;249;38;114mthen[0m
[38;2;248;248;242m                        tmp[0m[38;2;248;248;242m([0m[38;2;248;248;242mi[0m[38;2;248;248;242m)[0m[38;2;248;248;242m [0m[38;2;249;38;114m<=[0m[38;2;248;248;242m [0m[38;2;249;38;114mnot[0m[38;2;248;248;242m tmp[0m[38;2;248;248;242m([0m[38;2;248;248;242mi[0m[38;2;248;248;242m)[0m[38;2;248;248;242m;[0m
[38;2;248;248;242m                        i [0m[38;2;249;38;114m:=[0m[38;2;248;248;242m i [0m[38;2;249;38;114m+[0m[38;2;248;248;242m [0m[38;2;190;132;255m1[0m[38;2;248;248;242m;[0m
[38;2;248;248;242m                    [0m[38;2;249;38;114melse[0m
[38;2;248;248;242m                        state [0m[38;2;249;38;114m<=[0m[38;2;248;248;242m DONE[0m[38;2;248;248;242m;[0m
[38;2;248;248;242m                    [0m[38;2;249;38;114mend[0m[38;2;248;248;242m [0m[38;2;249;38;114mif[0m[38;2;248;248;242m;[0m

[38;2;248;248;242m                [0m[38;2;249;38;114mwhen[0m[38;2;248;248;242m DONE [0m[38;2;249;38;114m=>[0m
[38;2;248;248;242m                    flag [0m[38;2;249;38;114m<=[0m[38;2;248;248;242m [0m[38;2;190;132;255m'1'[0m[38;2;248;248;242m;[0m
[38;2;248;248;242m                    state [0m[38;2;249;38;114m<=[0m[38;2;248;248;242m IDLE[0m[38;2;248;248;242m;[0m

[38;2;248;248;242m                [0m[38;2;249;38;114mwhen[0m[38;2;248;248;242m [0m[38;2;249;38;114mothers[0m[38;2;248;248;242m [0m[38;2;249;38;114m=>[0m
[38;2;248;248;242m                    state [0m[38;2;249;38;114m<=[0m[38;2;248;248;242m IDLE[0m[38;2;248;248;242m;[0m
[38;2;248;248;242m            [0m[38;2;249;38;114mend[0m[38;2;248;248;242m [0m[38;2;249;38;114mcase[0m[38;2;248;248;242m;[0m
[38;2;248;248;242m        [0m[38;2;249;38;114mend[0m[38;2;248;248;242m [0m[38;2;249;38;114mif[0m[38;2;248;248;242m;[0m
[38;2;248;248;242m    [0m[38;2;249;38;114mend[0m[38;2;249;38;114m process[0m[38;2;248;248;242m;[0m

[38;2;248;248;242m    result [0m[38;2;249;38;114m<=[0m[38;2;248;248;242m tmp[0m[38;2;248;248;242m;[0m

[38;2;249;38;114mend[0m[38;2;248;248;242m [0m[38;2;166;226;46mBehavioral[0m[38;2;248;248;242m;[0m